//=======================================================
//  Module description
//=======================================================
`include "system_include.v"

module XXXX(

	//////////// CLOCK //////////
	input XXX,

	//  Only included if we're running with ModelSim
	`ifdef UNDER_TEST
		// Async reset
		input YYY,
	`endif
	
	//////////// LED //////////
	output ZZZ
);

//=======================================================
//  REG/WIRE declarations
//=======================================================

//=======================================================
//  Outputs
//=======================================================

//=======================================================
//  Structural coding
//=======================================================

//=======================================================
//  Procedural coding
//=======================================================
	
endmodule
